--ftp://www.cs.uregina.ca/pub/class/301/multiplexer/lecture.html
